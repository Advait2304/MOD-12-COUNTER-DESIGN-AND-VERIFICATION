package counter_pkg;
int no_of_transaction=1;
`include "transaction.sv"
`include "scoreboard.sv"
`include "driver.sv"
`include "generator.sv"
`include "wr_mon.sv"
`include "reference.sv"
`include "env.sv"
`include "test.sv"
`include "read_monitor.sv"
endpackage